`define BYTE 8
