module ex_t
(
    input logic clk_i,
    input logic rstn_i,

    input alu_op_t alu_op_i,
    output [(2*`BYTE)-1:0] alu_res_o
);


endmodule : ex_t
