module ex_t
(
    input logic clk_i,
    input logic rstn_i,

);


endmodule : ex_t
