module cpu_t
(
    input logic clk_i,
    input logic rstn_i

);

endmodule : cpu_t
