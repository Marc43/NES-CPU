package nes_cpu_pkg;
   
    int MEM_ADDR_SIZE = 16;         // 16 bits to index memory
    int BOOT_ADDR = 0;              // TODO Not really  
    int INSTR_SIZE_IN_BYTES = 16;   // So far 

endpackage : nes_cpu_pkg
