package nes_cpu_pkg;
   
    parameter int MEM_ADDR_SIZE = 16;         // 16 bits to index memory
    parameter int BOOT_ADDR = 0;              // TODO Not really  
    parameter int INSTR_SIZE_IN_BYTES = 2;    // So far 

endpackage : nes_cpu_pkg
